/* #### FONT0 #### */
reg [11:0] font0 [1709:0];

initial begin
font0[0] = 12'b000000000000;
font0[1] = 12'b000000000000;
font0[2] = 12'b000000000000;
font0[3] = 12'b000000000000;
font0[4] = 12'b000000000000;
font0[5] = 12'b000000000000;
font0[6] = 12'b000000000000;
font0[7] = 12'b000000000000;
font0[8] = 12'b000000000000;
font0[9] = 12'b000000000000;
font0[10] = 12'b000000000000;
font0[11] = 12'b000000000000;
font0[12] = 12'b000000000000;
font0[13] = 12'b000000000000;
font0[14] = 12'b000000000000;
font0[15] = 12'b000000000000;
font0[16] = 12'b000000000000;
font0[17] = 12'b000000000000;
font0[18] = 12'b000001000000;
font0[19] = 12'b000001000000;
font0[20] = 12'b000001000000;
font0[21] = 12'b000001100000;
font0[22] = 12'b000001100000;
font0[23] = 12'b000001100000;
font0[24] = 12'b000000000000;
font0[25] = 12'b000001100000;
font0[26] = 12'b000000000000;
font0[27] = 12'b000000000000;
font0[28] = 12'b000000000000;
font0[29] = 12'b000000000000;
font0[30] = 12'b000000000000;
font0[31] = 12'b000000000000;
font0[32] = 12'b000000000000;
font0[33] = 12'b000000000000;
font0[34] = 12'b000000000000;
font0[35] = 12'b000000000000;
font0[36] = 12'b000010100000;
font0[37] = 12'b000010100000;
font0[38] = 12'b000010100000;
font0[39] = 12'b000000000000;
font0[40] = 12'b000000000000;
font0[41] = 12'b000000000000;
font0[42] = 12'b000000000000;
font0[43] = 12'b000000000000;
font0[44] = 12'b000000000000;
font0[45] = 12'b000000000000;
font0[46] = 12'b000000000000;
font0[47] = 12'b000000000000;
font0[48] = 12'b000000000000;
font0[49] = 12'b000000000000;
font0[50] = 12'b000000000000;
font0[51] = 12'b000000000000;
font0[52] = 12'b000000000000;
font0[53] = 12'b000000000000;
font0[54] = 12'b000100010000;
font0[55] = 12'b000100010000;
font0[56] = 12'b001111111100;
font0[57] = 12'b000100010000;
font0[58] = 12'b000110011000;
font0[59] = 12'b001111111100;
font0[60] = 12'b000110011000;
font0[61] = 12'b000110011000;
font0[62] = 12'b000000000000;
font0[63] = 12'b000000000000;
font0[64] = 12'b000000000000;
font0[65] = 12'b000000000000;
font0[66] = 12'b000000000000;
font0[67] = 12'b000000000000;
font0[68] = 12'b000000000000;
font0[69] = 12'b000000000000;
font0[70] = 12'b000000000000;
font0[71] = 12'b000000000000;
font0[72] = 12'b000011111000;
font0[73] = 12'b000100100000;
font0[74] = 12'b000100100000;
font0[75] = 12'b000100100000;
font0[76] = 12'b000011111000;
font0[77] = 12'b000000111000;
font0[78] = 12'b000000111000;
font0[79] = 12'b000111111000;
font0[80] = 12'b000000100000;
font0[81] = 12'b000000000000;
font0[82] = 12'b000000000000;
font0[83] = 12'b000000000000;
font0[84] = 12'b000000000000;
font0[85] = 12'b000000000000;
font0[86] = 12'b000000000000;
font0[87] = 12'b000000000000;
font0[88] = 12'b000000000000;
font0[89] = 12'b000000000000;
font0[90] = 12'b001110000000;
font0[91] = 12'b001010100000;
font0[92] = 12'b001111100000;
font0[93] = 12'b000001000000;
font0[94] = 12'b000011000000;
font0[95] = 12'b000011011100;
font0[96] = 12'b000110011100;
font0[97] = 12'b000110011100;
font0[98] = 12'b000000000000;
font0[99] = 12'b000000000000;
font0[100] = 12'b000000000000;
font0[101] = 12'b000000000000;
font0[102] = 12'b000000000000;
font0[103] = 12'b000000000000;
font0[104] = 12'b000000000000;
font0[105] = 12'b000000000000;
font0[106] = 12'b000000000000;
font0[107] = 12'b000000000000;
font0[108] = 12'b000111100000;
font0[109] = 12'b001000010000;
font0[110] = 12'b001000010000;
font0[111] = 12'b001000010000;
font0[112] = 12'b001111111000;
font0[113] = 12'b001100010000;
font0[114] = 12'b001100010000;
font0[115] = 12'b000111111100;
font0[116] = 12'b000000000000;
font0[117] = 12'b000000000000;
font0[118] = 12'b000000000000;
font0[119] = 12'b000000000000;
font0[120] = 12'b000000000000;
font0[121] = 12'b000000000000;
font0[122] = 12'b000000000000;
font0[123] = 12'b000000000000;
font0[124] = 12'b000000000000;
font0[125] = 12'b000000000000;
font0[126] = 12'b000001000000;
font0[127] = 12'b000001000000;
font0[128] = 12'b000001000000;
font0[129] = 12'b000000000000;
font0[130] = 12'b000000000000;
font0[131] = 12'b000000000000;
font0[132] = 12'b000000000000;
font0[133] = 12'b000000000000;
font0[134] = 12'b000000000000;
font0[135] = 12'b000000000000;
font0[136] = 12'b000000000000;
font0[137] = 12'b000000000000;
font0[138] = 12'b000000000000;
font0[139] = 12'b000000000000;
font0[140] = 12'b000000000000;
font0[141] = 12'b000000000000;
font0[142] = 12'b000000000000;
font0[143] = 12'b000000000000;
font0[144] = 12'b000001110000;
font0[145] = 12'b000010000000;
font0[146] = 12'b000010000000;
font0[147] = 12'b000011000000;
font0[148] = 12'b000011000000;
font0[149] = 12'b000011000000;
font0[150] = 12'b000011000000;
font0[151] = 12'b000001110000;
font0[152] = 12'b000000000000;
font0[153] = 12'b000000000000;
font0[154] = 12'b000000000000;
font0[155] = 12'b000000000000;
font0[156] = 12'b000000000000;
font0[157] = 12'b000000000000;
font0[158] = 12'b000000000000;
font0[159] = 12'b000000000000;
font0[160] = 12'b000000000000;
font0[161] = 12'b000000000000;
font0[162] = 12'b000011100000;
font0[163] = 12'b000000010000;
font0[164] = 12'b000000010000;
font0[165] = 12'b000000110000;
font0[166] = 12'b000000110000;
font0[167] = 12'b000000110000;
font0[168] = 12'b000000110000;
font0[169] = 12'b000011100000;
font0[170] = 12'b000000000000;
font0[171] = 12'b000000000000;
font0[172] = 12'b000000000000;
font0[173] = 12'b000000000000;
font0[174] = 12'b000000000000;
font0[175] = 12'b000000000000;
font0[176] = 12'b000000000000;
font0[177] = 12'b000000000000;
font0[178] = 12'b000000000000;
font0[179] = 12'b000000000000;
font0[180] = 12'b000000000000;
font0[181] = 12'b000000000000;
font0[182] = 12'b000111100000;
font0[183] = 12'b000011000000;
font0[184] = 12'b000111110000;
font0[185] = 12'b000111100000;
font0[186] = 12'b000000000000;
font0[187] = 12'b000000000000;
font0[188] = 12'b000000000000;
font0[189] = 12'b000000000000;
font0[190] = 12'b000000000000;
font0[191] = 12'b000000000000;
font0[192] = 12'b000000000000;
font0[193] = 12'b000000000000;
font0[194] = 12'b000000000000;
font0[195] = 12'b000000000000;
font0[196] = 12'b000000000000;
font0[197] = 12'b000000000000;
font0[198] = 12'b000000000000;
font0[199] = 12'b000001000000;
font0[200] = 12'b000001000000;
font0[201] = 12'b000001000000;
font0[202] = 12'b001111111000;
font0[203] = 12'b000001100000;
font0[204] = 12'b000001100000;
font0[205] = 12'b000001100000;
font0[206] = 12'b000000000000;
font0[207] = 12'b000000000000;
font0[208] = 12'b000000000000;
font0[209] = 12'b000000000000;
font0[210] = 12'b000000000000;
font0[211] = 12'b000000000000;
font0[212] = 12'b000000000000;
font0[213] = 12'b000000000000;
font0[214] = 12'b000000000000;
font0[215] = 12'b000000000000;
font0[216] = 12'b000000000000;
font0[217] = 12'b000000000000;
font0[218] = 12'b000000000000;
font0[219] = 12'b000000000000;
font0[220] = 12'b000000000000;
font0[221] = 12'b000000000000;
font0[222] = 12'b000000000000;
font0[223] = 12'b000001100000;
font0[224] = 12'b000000100000;
font0[225] = 12'b000000100000;
font0[226] = 12'b000000000000;
font0[227] = 12'b000000000000;
font0[228] = 12'b000000000000;
font0[229] = 12'b000000000000;
font0[230] = 12'b000000000000;
font0[231] = 12'b000000000000;
font0[232] = 12'b000000000000;
font0[233] = 12'b000000000000;
font0[234] = 12'b000000000000;
font0[235] = 12'b000000000000;
font0[236] = 12'b000000000000;
font0[237] = 12'b000000000000;
font0[238] = 12'b001111111000;
font0[239] = 12'b000000000000;
font0[240] = 12'b000000000000;
font0[241] = 12'b000000000000;
font0[242] = 12'b000000000000;
font0[243] = 12'b000000000000;
font0[244] = 12'b000000000000;
font0[245] = 12'b000000000000;
font0[246] = 12'b000000000000;
font0[247] = 12'b000000000000;
font0[248] = 12'b000000000000;
font0[249] = 12'b000000000000;
font0[250] = 12'b000000000000;
font0[251] = 12'b000000000000;
font0[252] = 12'b000000000000;
font0[253] = 12'b000000000000;
font0[254] = 12'b000000000000;
font0[255] = 12'b000000000000;
font0[256] = 12'b000000000000;
font0[257] = 12'b000000000000;
font0[258] = 12'b000000000000;
font0[259] = 12'b000001100000;
font0[260] = 12'b000000000000;
font0[261] = 12'b000000000000;
font0[262] = 12'b000000000000;
font0[263] = 12'b000000000000;
font0[264] = 12'b000000000000;
font0[265] = 12'b000000000000;
font0[266] = 12'b000000000000;
font0[267] = 12'b000000000000;
font0[268] = 12'b000000000000;
font0[269] = 12'b000000000000;
font0[270] = 12'b000000000000;
font0[271] = 12'b000000010000;
font0[272] = 12'b000000010000;
font0[273] = 12'b000000100000;
font0[274] = 12'b000001100000;
font0[275] = 12'b000001100000;
font0[276] = 12'b000011000000;
font0[277] = 12'b000011000000;
font0[278] = 12'b000000000000;
font0[279] = 12'b000000000000;
font0[280] = 12'b000000000000;
font0[281] = 12'b000000000000;
font0[282] = 12'b000000000000;
font0[283] = 12'b000000000000;
font0[284] = 12'b000000000000;
font0[285] = 12'b000000000000;
font0[286] = 12'b000000000000;
font0[287] = 12'b000000000000;
font0[288] = 12'b000011110000;
font0[289] = 12'b000100011000;
font0[290] = 12'b000100011000;
font0[291] = 12'b000110011000;
font0[292] = 12'b000110011000;
font0[293] = 12'b000110001000;
font0[294] = 12'b000110001000;
font0[295] = 12'b000011110000;
font0[296] = 12'b000000000000;
font0[297] = 12'b000000000000;
font0[298] = 12'b000000000000;
font0[299] = 12'b000000000000;
font0[300] = 12'b000000000000;
font0[301] = 12'b000000000000;
font0[302] = 12'b000000000000;
font0[303] = 12'b000000000000;
font0[304] = 12'b000000000000;
font0[305] = 12'b000000000000;
font0[306] = 12'b000011100000;
font0[307] = 12'b000000100000;
font0[308] = 12'b000000100000;
font0[309] = 12'b000001100000;
font0[310] = 12'b000001100000;
font0[311] = 12'b000001100000;
font0[312] = 12'b000001100000;
font0[313] = 12'b000111111000;
font0[314] = 12'b000000000000;
font0[315] = 12'b000000000000;
font0[316] = 12'b000000000000;
font0[317] = 12'b000000000000;
font0[318] = 12'b000000000000;
font0[319] = 12'b000000000000;
font0[320] = 12'b000000000000;
font0[321] = 12'b000000000000;
font0[322] = 12'b000000000000;
font0[323] = 12'b000000000000;
font0[324] = 12'b000111110000;
font0[325] = 12'b000000001000;
font0[326] = 12'b000000001000;
font0[327] = 12'b000000001000;
font0[328] = 12'b000111110000;
font0[329] = 12'b000110000000;
font0[330] = 12'b000110000000;
font0[331] = 12'b000111111000;
font0[332] = 12'b000000000000;
font0[333] = 12'b000000000000;
font0[334] = 12'b000000000000;
font0[335] = 12'b000000000000;
font0[336] = 12'b000000000000;
font0[337] = 12'b000000000000;
font0[338] = 12'b000000000000;
font0[339] = 12'b000000000000;
font0[340] = 12'b000000000000;
font0[341] = 12'b000000000000;
font0[342] = 12'b001111110000;
font0[343] = 12'b000000001000;
font0[344] = 12'b000000001000;
font0[345] = 12'b000000001000;
font0[346] = 12'b000011111000;
font0[347] = 12'b000000011000;
font0[348] = 12'b000000011000;
font0[349] = 12'b001111110000;
font0[350] = 12'b000000000000;
font0[351] = 12'b000000000000;
font0[352] = 12'b000000000000;
font0[353] = 12'b000000000000;
font0[354] = 12'b000000000000;
font0[355] = 12'b000000000000;
font0[356] = 12'b000000000000;
font0[357] = 12'b000000000000;
font0[358] = 12'b000000000000;
font0[359] = 12'b000000000000;
font0[360] = 12'b000100001000;
font0[361] = 12'b000100001000;
font0[362] = 12'b000100001000;
font0[363] = 12'b000100001000;
font0[364] = 12'b000111111000;
font0[365] = 12'b000000011000;
font0[366] = 12'b000000011000;
font0[367] = 12'b000000011000;
font0[368] = 12'b000000000000;
font0[369] = 12'b000000000000;
font0[370] = 12'b000000000000;
font0[371] = 12'b000000000000;
font0[372] = 12'b000000000000;
font0[373] = 12'b000000000000;
font0[374] = 12'b000000000000;
font0[375] = 12'b000000000000;
font0[376] = 12'b000000000000;
font0[377] = 12'b000000000000;
font0[378] = 12'b000111111000;
font0[379] = 12'b000100000000;
font0[380] = 12'b000100000000;
font0[381] = 12'b000100000000;
font0[382] = 12'b000111111000;
font0[383] = 12'b000000011000;
font0[384] = 12'b000000011000;
font0[385] = 12'b000111111000;
font0[386] = 12'b000000000000;
font0[387] = 12'b000000000000;
font0[388] = 12'b000000000000;
font0[389] = 12'b000000000000;
font0[390] = 12'b000000000000;
font0[391] = 12'b000000000000;
font0[392] = 12'b000000000000;
font0[393] = 12'b000000000000;
font0[394] = 12'b000000000000;
font0[395] = 12'b000000000000;
font0[396] = 12'b000011110000;
font0[397] = 12'b000100000000;
font0[398] = 12'b000100000000;
font0[399] = 12'b000100000000;
font0[400] = 12'b000111111000;
font0[401] = 12'b000110001000;
font0[402] = 12'b000110001000;
font0[403] = 12'b000011110000;
font0[404] = 12'b000000000000;
font0[405] = 12'b000000000000;
font0[406] = 12'b000000000000;
font0[407] = 12'b000000000000;
font0[408] = 12'b000000000000;
font0[409] = 12'b000000000000;
font0[410] = 12'b000000000000;
font0[411] = 12'b000000000000;
font0[412] = 12'b000000000000;
font0[413] = 12'b000000000000;
font0[414] = 12'b001111111000;
font0[415] = 12'b000000001000;
font0[416] = 12'b000000001000;
font0[417] = 12'b000000001000;
font0[418] = 12'b000000011000;
font0[419] = 12'b000000011000;
font0[420] = 12'b000000011000;
font0[421] = 12'b000000011000;
font0[422] = 12'b000000000000;
font0[423] = 12'b000000000000;
font0[424] = 12'b000000000000;
font0[425] = 12'b000000000000;
font0[426] = 12'b000000000000;
font0[427] = 12'b000000000000;
font0[428] = 12'b000000000000;
font0[429] = 12'b000000000000;
font0[430] = 12'b000000000000;
font0[431] = 12'b000000000000;
font0[432] = 12'b000011111000;
font0[433] = 12'b000100001000;
font0[434] = 12'b000100001000;
font0[435] = 12'b000100001000;
font0[436] = 12'b000111111000;
font0[437] = 12'b000110011000;
font0[438] = 12'b000110011000;
font0[439] = 12'b000011111000;
font0[440] = 12'b000000000000;
font0[441] = 12'b000000000000;
font0[442] = 12'b000000000000;
font0[443] = 12'b000000000000;
font0[444] = 12'b000000000000;
font0[445] = 12'b000000000000;
font0[446] = 12'b000000000000;
font0[447] = 12'b000000000000;
font0[448] = 12'b000000000000;
font0[449] = 12'b000000000000;
font0[450] = 12'b000011110000;
font0[451] = 12'b000100001000;
font0[452] = 12'b000100001000;
font0[453] = 12'b000100001000;
font0[454] = 12'b000011111000;
font0[455] = 12'b000000011000;
font0[456] = 12'b000000011000;
font0[457] = 12'b000011110000;
font0[458] = 12'b000000000000;
font0[459] = 12'b000000000000;
font0[460] = 12'b000000000000;
font0[461] = 12'b000000000000;
font0[462] = 12'b000000000000;
font0[463] = 12'b000000000000;
font0[464] = 12'b000000000000;
font0[465] = 12'b000000000000;
font0[466] = 12'b000000000000;
font0[467] = 12'b000000000000;
font0[468] = 12'b000000000000;
font0[469] = 12'b000000000000;
font0[470] = 12'b000001100000;
font0[471] = 12'b000000000000;
font0[472] = 12'b000000000000;
font0[473] = 12'b000001100000;
font0[474] = 12'b000000000000;
font0[475] = 12'b000000000000;
font0[476] = 12'b000000000000;
font0[477] = 12'b000000000000;
font0[478] = 12'b000000000000;
font0[479] = 12'b000000000000;
font0[480] = 12'b000000000000;
font0[481] = 12'b000000000000;
font0[482] = 12'b000000000000;
font0[483] = 12'b000000000000;
font0[484] = 12'b000000000000;
font0[485] = 12'b000000000000;
font0[486] = 12'b000000000000;
font0[487] = 12'b000000000000;
font0[488] = 12'b000001100000;
font0[489] = 12'b000000000000;
font0[490] = 12'b000000000000;
font0[491] = 12'b000000000000;
font0[492] = 12'b000000000000;
font0[493] = 12'b000001100000;
font0[494] = 12'b000000100000;
font0[495] = 12'b000000100000;
font0[496] = 12'b000000000000;
font0[497] = 12'b000000000000;
font0[498] = 12'b000000000000;
font0[499] = 12'b000000000000;
font0[500] = 12'b000000000000;
font0[501] = 12'b000000000000;
font0[502] = 12'b000000000000;
font0[503] = 12'b000000000000;
font0[504] = 12'b000000000000;
font0[505] = 12'b000000010000;
font0[506] = 12'b000000100000;
font0[507] = 12'b000001000000;
font0[508] = 12'b000001100000;
font0[509] = 12'b000001110000;
font0[510] = 12'b000000010000;
font0[511] = 12'b000000000000;
font0[512] = 12'b000000000000;
font0[513] = 12'b000000000000;
font0[514] = 12'b000000000000;
font0[515] = 12'b000000000000;
font0[516] = 12'b000000000000;
font0[517] = 12'b000000000000;
font0[518] = 12'b000000000000;
font0[519] = 12'b000000000000;
font0[520] = 12'b000000000000;
font0[521] = 12'b000000000000;
font0[522] = 12'b000000000000;
font0[523] = 12'b000000000000;
font0[524] = 12'b001111111000;
font0[525] = 12'b000000000000;
font0[526] = 12'b000000000000;
font0[527] = 12'b001111111000;
font0[528] = 12'b000000000000;
font0[529] = 12'b000000000000;
font0[530] = 12'b000000000000;
font0[531] = 12'b000000000000;
font0[532] = 12'b000000000000;
font0[533] = 12'b000000000000;
font0[534] = 12'b000000000000;
font0[535] = 12'b000000000000;
font0[536] = 12'b000000000000;
font0[537] = 12'b000000000000;
font0[538] = 12'b000000000000;
font0[539] = 12'b000000000000;
font0[540] = 12'b000000000000;
font0[541] = 12'b000010000000;
font0[542] = 12'b000001000000;
font0[543] = 12'b000000100000;
font0[544] = 12'b000001100000;
font0[545] = 12'b000011100000;
font0[546] = 12'b000010000000;
font0[547] = 12'b000000000000;
font0[548] = 12'b000000000000;
font0[549] = 12'b000000000000;
font0[550] = 12'b000000000000;
font0[551] = 12'b000000000000;
font0[552] = 12'b000000000000;
font0[553] = 12'b000000000000;
font0[554] = 12'b000000000000;
font0[555] = 12'b000000000000;
font0[556] = 12'b000000000000;
font0[557] = 12'b000000000000;
font0[558] = 12'b000111110000;
font0[559] = 12'b001100001000;
font0[560] = 12'b000000001000;
font0[561] = 12'b000000001000;
font0[562] = 12'b000001110000;
font0[563] = 12'b000001100000;
font0[564] = 12'b000001100000;
font0[565] = 12'b000001100000;
font0[566] = 12'b000000000000;
font0[567] = 12'b000000000000;
font0[568] = 12'b000000000000;
font0[569] = 12'b000000000000;
font0[570] = 12'b000000000000;
font0[571] = 12'b000000000000;
font0[572] = 12'b000000000000;
font0[573] = 12'b000000000000;
font0[574] = 12'b000000000000;
font0[575] = 12'b000000000000;
font0[576] = 12'b000111111000;
font0[577] = 12'b000100001000;
font0[578] = 12'b000101111000;
font0[579] = 12'b000111111000;
font0[580] = 12'b000111111000;
font0[581] = 12'b000111111000;
font0[582] = 12'b000110000000;
font0[583] = 12'b000111110000;
font0[584] = 12'b000000000000;
font0[585] = 12'b000000000000;
font0[586] = 12'b000000000000;
font0[587] = 12'b000000000000;
font0[588] = 12'b000000000000;
font0[589] = 12'b000000000000;
font0[590] = 12'b000000000000;
font0[591] = 12'b000000000000;
font0[592] = 12'b000000000000;
font0[593] = 12'b000000000000;
font0[594] = 12'b000111111000;
font0[595] = 12'b000100001000;
font0[596] = 12'b000100001000;
font0[597] = 12'b000100001000;
font0[598] = 12'b000111111000;
font0[599] = 12'b000110011000;
font0[600] = 12'b000110011000;
font0[601] = 12'b000110011000;
font0[602] = 12'b000000000000;
font0[603] = 12'b000000000000;
font0[604] = 12'b000000000000;
font0[605] = 12'b000000000000;
font0[606] = 12'b000000000000;
font0[607] = 12'b000000000000;
font0[608] = 12'b000000000000;
font0[609] = 12'b000000000000;
font0[610] = 12'b000000000000;
font0[611] = 12'b000000000000;
font0[612] = 12'b000111110000;
font0[613] = 12'b000100001000;
font0[614] = 12'b000100001000;
font0[615] = 12'b000100001000;
font0[616] = 12'b000111111000;
font0[617] = 12'b000110001000;
font0[618] = 12'b000110001000;
font0[619] = 12'b000111110000;
font0[620] = 12'b000000000000;
font0[621] = 12'b000000000000;
font0[622] = 12'b000000000000;
font0[623] = 12'b000000000000;
font0[624] = 12'b000000000000;
font0[625] = 12'b000000000000;
font0[626] = 12'b000000000000;
font0[627] = 12'b000000000000;
font0[628] = 12'b000000000000;
font0[629] = 12'b000000000000;
font0[630] = 12'b000111111000;
font0[631] = 12'b001000000000;
font0[632] = 12'b001000000000;
font0[633] = 12'b001100000000;
font0[634] = 12'b001100000000;
font0[635] = 12'b001100000000;
font0[636] = 12'b001100000000;
font0[637] = 12'b000111111000;
font0[638] = 12'b000000000000;
font0[639] = 12'b000000000000;
font0[640] = 12'b000000000000;
font0[641] = 12'b000000000000;
font0[642] = 12'b000000000000;
font0[643] = 12'b000000000000;
font0[644] = 12'b000000000000;
font0[645] = 12'b000000000000;
font0[646] = 12'b000000000000;
font0[647] = 12'b000000000000;
font0[648] = 12'b000111110000;
font0[649] = 12'b000100001000;
font0[650] = 12'b000100001000;
font0[651] = 12'b000110001000;
font0[652] = 12'b000110001000;
font0[653] = 12'b000110001000;
font0[654] = 12'b000110001000;
font0[655] = 12'b000111110000;
font0[656] = 12'b000000000000;
font0[657] = 12'b000000000000;
font0[658] = 12'b000000000000;
font0[659] = 12'b000000000000;
font0[660] = 12'b000000000000;
font0[661] = 12'b000000000000;
font0[662] = 12'b000000000000;
font0[663] = 12'b000000000000;
font0[664] = 12'b000000000000;
font0[665] = 12'b000000000000;
font0[666] = 12'b001111111000;
font0[667] = 12'b001000000000;
font0[668] = 12'b001000000000;
font0[669] = 12'b001000000000;
font0[670] = 12'b001111110000;
font0[671] = 12'b001100000000;
font0[672] = 12'b001100000000;
font0[673] = 12'b001111111000;
font0[674] = 12'b000000000000;
font0[675] = 12'b000000000000;
font0[676] = 12'b000000000000;
font0[677] = 12'b000000000000;
font0[678] = 12'b000000000000;
font0[679] = 12'b000000000000;
font0[680] = 12'b000000000000;
font0[681] = 12'b000000000000;
font0[682] = 12'b000000000000;
font0[683] = 12'b000000000000;
font0[684] = 12'b001111111000;
font0[685] = 12'b001000000000;
font0[686] = 12'b001000000000;
font0[687] = 12'b001000000000;
font0[688] = 12'b001111110000;
font0[689] = 12'b001100000000;
font0[690] = 12'b001100000000;
font0[691] = 12'b001100000000;
font0[692] = 12'b000000000000;
font0[693] = 12'b000000000000;
font0[694] = 12'b000000000000;
font0[695] = 12'b000000000000;
font0[696] = 12'b000000000000;
font0[697] = 12'b000000000000;
font0[698] = 12'b000000000000;
font0[699] = 12'b000000000000;
font0[700] = 12'b000000000000;
font0[701] = 12'b000000000000;
font0[702] = 12'b000011110000;
font0[703] = 12'b000100000000;
font0[704] = 12'b000100000000;
font0[705] = 12'b000100000000;
font0[706] = 12'b000110111000;
font0[707] = 12'b000110001000;
font0[708] = 12'b000110001000;
font0[709] = 12'b000011110000;
font0[710] = 12'b000000000000;
font0[711] = 12'b000000000000;
font0[712] = 12'b000000000000;
font0[713] = 12'b000000000000;
font0[714] = 12'b000000000000;
font0[715] = 12'b000000000000;
font0[716] = 12'b000000000000;
font0[717] = 12'b000000000000;
font0[718] = 12'b000000000000;
font0[719] = 12'b000000000000;
font0[720] = 12'b000100001000;
font0[721] = 12'b000100001000;
font0[722] = 12'b000100001000;
font0[723] = 12'b000100001000;
font0[724] = 12'b000111111000;
font0[725] = 12'b000110011000;
font0[726] = 12'b000110011000;
font0[727] = 12'b000110011000;
font0[728] = 12'b000000000000;
font0[729] = 12'b000000000000;
font0[730] = 12'b000000000000;
font0[731] = 12'b000000000000;
font0[732] = 12'b000000000000;
font0[733] = 12'b000000000000;
font0[734] = 12'b000000000000;
font0[735] = 12'b000000000000;
font0[736] = 12'b000000000000;
font0[737] = 12'b000000000000;
font0[738] = 12'b000011110000;
font0[739] = 12'b000000100000;
font0[740] = 12'b000000100000;
font0[741] = 12'b000001100000;
font0[742] = 12'b000001100000;
font0[743] = 12'b000001100000;
font0[744] = 12'b000001100000;
font0[745] = 12'b000011110000;
font0[746] = 12'b000000000000;
font0[747] = 12'b000000000000;
font0[748] = 12'b000000000000;
font0[749] = 12'b000000000000;
font0[750] = 12'b000000000000;
font0[751] = 12'b000000000000;
font0[752] = 12'b000000000000;
font0[753] = 12'b000000000000;
font0[754] = 12'b000000000000;
font0[755] = 12'b000000000000;
font0[756] = 12'b000111111000;
font0[757] = 12'b000000001000;
font0[758] = 12'b000000001000;
font0[759] = 12'b000000011000;
font0[760] = 12'b000100011000;
font0[761] = 12'b000100011000;
font0[762] = 12'b000100011000;
font0[763] = 12'b000011110000;
font0[764] = 12'b000000000000;
font0[765] = 12'b000000000000;
font0[766] = 12'b000000000000;
font0[767] = 12'b000000000000;
font0[768] = 12'b000000000000;
font0[769] = 12'b000000000000;
font0[770] = 12'b000000000000;
font0[771] = 12'b000000000000;
font0[772] = 12'b000000000000;
font0[773] = 12'b000000000000;
font0[774] = 12'b000100001000;
font0[775] = 12'b000100001000;
font0[776] = 12'b000100010000;
font0[777] = 12'b000100110000;
font0[778] = 12'b000110110000;
font0[779] = 12'b000110010000;
font0[780] = 12'b000110001000;
font0[781] = 12'b000110001000;
font0[782] = 12'b000000000000;
font0[783] = 12'b000000000000;
font0[784] = 12'b000000000000;
font0[785] = 12'b000000000000;
font0[786] = 12'b000000000000;
font0[787] = 12'b000000000000;
font0[788] = 12'b000000000000;
font0[789] = 12'b000000000000;
font0[790] = 12'b000000000000;
font0[791] = 12'b000000000000;
font0[792] = 12'b001000000000;
font0[793] = 12'b001000000000;
font0[794] = 12'b001000000000;
font0[795] = 12'b001100000000;
font0[796] = 12'b001100000000;
font0[797] = 12'b001100000000;
font0[798] = 12'b001100000000;
font0[799] = 12'b001111111000;
font0[800] = 12'b000000000000;
font0[801] = 12'b000000000000;
font0[802] = 12'b000000000000;
font0[803] = 12'b000000000000;
font0[804] = 12'b000000000000;
font0[805] = 12'b000000000000;
font0[806] = 12'b000000000000;
font0[807] = 12'b000000000000;
font0[808] = 12'b000000000000;
font0[809] = 12'b000000000000;
font0[810] = 12'b000100001000;
font0[811] = 12'b000100001000;
font0[812] = 12'b000100001000;
font0[813] = 12'b000110011000;
font0[814] = 12'b000111111000;
font0[815] = 12'b000110111000;
font0[816] = 12'b000110011000;
font0[817] = 12'b000110011000;
font0[818] = 12'b000000000000;
font0[819] = 12'b000000000000;
font0[820] = 12'b000000000000;
font0[821] = 12'b000000000000;
font0[822] = 12'b000000000000;
font0[823] = 12'b000000000000;
font0[824] = 12'b000000000000;
font0[825] = 12'b000000000000;
font0[826] = 12'b000000000000;
font0[827] = 12'b000000000000;
font0[828] = 12'b000100001000;
font0[829] = 12'b000100001000;
font0[830] = 12'b000110001000;
font0[831] = 12'b000111001000;
font0[832] = 12'b000110111000;
font0[833] = 12'b000110011000;
font0[834] = 12'b000110001000;
font0[835] = 12'b000110001000;
font0[836] = 12'b000000000000;
font0[837] = 12'b000000000000;
font0[838] = 12'b000000000000;
font0[839] = 12'b000000000000;
font0[840] = 12'b000000000000;
font0[841] = 12'b000000000000;
font0[842] = 12'b000000000000;
font0[843] = 12'b000000000000;
font0[844] = 12'b000000000000;
font0[845] = 12'b000000000000;
font0[846] = 12'b000011110000;
font0[847] = 12'b000100001000;
font0[848] = 12'b000100001000;
font0[849] = 12'b000110011000;
font0[850] = 12'b000110011000;
font0[851] = 12'b000110011000;
font0[852] = 12'b000110011000;
font0[853] = 12'b000011110000;
font0[854] = 12'b000000000000;
font0[855] = 12'b000000000000;
font0[856] = 12'b000000000000;
font0[857] = 12'b000000000000;
font0[858] = 12'b000000000000;
font0[859] = 12'b000000000000;
font0[860] = 12'b000000000000;
font0[861] = 12'b000000000000;
font0[862] = 12'b000000000000;
font0[863] = 12'b000000000000;
font0[864] = 12'b000111110000;
font0[865] = 12'b000100001000;
font0[866] = 12'b000100001000;
font0[867] = 12'b000100001000;
font0[868] = 12'b000111110000;
font0[869] = 12'b000110000000;
font0[870] = 12'b000110000000;
font0[871] = 12'b000110000000;
font0[872] = 12'b000000000000;
font0[873] = 12'b000000000000;
font0[874] = 12'b000000000000;
font0[875] = 12'b000000000000;
font0[876] = 12'b000000000000;
font0[877] = 12'b000000000000;
font0[878] = 12'b000000000000;
font0[879] = 12'b000000000000;
font0[880] = 12'b000000000000;
font0[881] = 12'b000000000000;
font0[882] = 12'b000011110000;
font0[883] = 12'b000100001000;
font0[884] = 12'b000100001000;
font0[885] = 12'b000100011000;
font0[886] = 12'b000100011000;
font0[887] = 12'b000100011000;
font0[888] = 12'b000100011000;
font0[889] = 12'b000011111000;
font0[890] = 12'b000000000000;
font0[891] = 12'b000000000000;
font0[892] = 12'b000000000000;
font0[893] = 12'b000000000000;
font0[894] = 12'b000000000000;
font0[895] = 12'b000000000000;
font0[896] = 12'b000000000000;
font0[897] = 12'b000000000000;
font0[898] = 12'b000000000000;
font0[899] = 12'b000000000000;
font0[900] = 12'b000111110000;
font0[901] = 12'b000100001000;
font0[902] = 12'b000100001000;
font0[903] = 12'b000100001000;
font0[904] = 12'b000111110000;
font0[905] = 12'b000110010000;
font0[906] = 12'b000110001000;
font0[907] = 12'b000110001000;
font0[908] = 12'b000000000000;
font0[909] = 12'b000000000000;
font0[910] = 12'b000000000000;
font0[911] = 12'b000000000000;
font0[912] = 12'b000000000000;
font0[913] = 12'b000000000000;
font0[914] = 12'b000000000000;
font0[915] = 12'b000000000000;
font0[916] = 12'b000000000000;
font0[917] = 12'b000000000000;
font0[918] = 12'b000011111000;
font0[919] = 12'b000100000000;
font0[920] = 12'b000100000000;
font0[921] = 12'b000100000000;
font0[922] = 12'b000011111000;
font0[923] = 12'b000000011000;
font0[924] = 12'b000000011000;
font0[925] = 12'b000111111000;
font0[926] = 12'b000000000000;
font0[927] = 12'b000000000000;
font0[928] = 12'b000000000000;
font0[929] = 12'b000000000000;
font0[930] = 12'b000000000000;
font0[931] = 12'b000000000000;
font0[932] = 12'b000000000000;
font0[933] = 12'b000000000000;
font0[934] = 12'b000000000000;
font0[935] = 12'b000000000000;
font0[936] = 12'b001111111000;
font0[937] = 12'b000001000000;
font0[938] = 12'b000001000000;
font0[939] = 12'b000001000000;
font0[940] = 12'b000011000000;
font0[941] = 12'b000011000000;
font0[942] = 12'b000011000000;
font0[943] = 12'b000011000000;
font0[944] = 12'b000000000000;
font0[945] = 12'b000000000000;
font0[946] = 12'b000000000000;
font0[947] = 12'b000000000000;
font0[948] = 12'b000000000000;
font0[949] = 12'b000000000000;
font0[950] = 12'b000000000000;
font0[951] = 12'b000000000000;
font0[952] = 12'b000000000000;
font0[953] = 12'b000000000000;
font0[954] = 12'b000100001000;
font0[955] = 12'b000100001000;
font0[956] = 12'b000100001000;
font0[957] = 12'b000110011000;
font0[958] = 12'b000110011000;
font0[959] = 12'b000110011000;
font0[960] = 12'b000110011000;
font0[961] = 12'b000011110000;
font0[962] = 12'b000000000000;
font0[963] = 12'b000000000000;
font0[964] = 12'b000000000000;
font0[965] = 12'b000000000000;
font0[966] = 12'b000000000000;
font0[967] = 12'b000000000000;
font0[968] = 12'b000000000000;
font0[969] = 12'b000000000000;
font0[970] = 12'b000000000000;
font0[971] = 12'b000000000000;
font0[972] = 12'b000100001000;
font0[973] = 12'b000100001000;
font0[974] = 12'b000100001000;
font0[975] = 12'b000100001000;
font0[976] = 12'b000110011000;
font0[977] = 12'b000010010000;
font0[978] = 12'b000011110000;
font0[979] = 12'b000001100000;
font0[980] = 12'b000000000000;
font0[981] = 12'b000000000000;
font0[982] = 12'b000000000000;
font0[983] = 12'b000000000000;
font0[984] = 12'b000000000000;
font0[985] = 12'b000000000000;
font0[986] = 12'b000000000000;
font0[987] = 12'b000000000000;
font0[988] = 12'b000000000000;
font0[989] = 12'b000000000000;
font0[990] = 12'b000100001000;
font0[991] = 12'b000100001000;
font0[992] = 12'b000100101000;
font0[993] = 12'b000110111000;
font0[994] = 12'b000110111000;
font0[995] = 12'b000110111000;
font0[996] = 12'b000110111000;
font0[997] = 12'b000011110000;
font0[998] = 12'b000000000000;
font0[999] = 12'b000000000000;
font0[1000] = 12'b000000000000;
font0[1001] = 12'b000000000000;
font0[1002] = 12'b000000000000;
font0[1003] = 12'b000000000000;
font0[1004] = 12'b000000000000;
font0[1005] = 12'b000000000000;
font0[1006] = 12'b000000000000;
font0[1007] = 12'b000000000000;
font0[1008] = 12'b000100001000;
font0[1009] = 12'b000100001000;
font0[1010] = 12'b000010010000;
font0[1011] = 12'b000011110000;
font0[1012] = 12'b000011110000;
font0[1013] = 12'b000010010000;
font0[1014] = 12'b000110011000;
font0[1015] = 12'b000110011000;
font0[1016] = 12'b000000000000;
font0[1017] = 12'b000000000000;
font0[1018] = 12'b000000000000;
font0[1019] = 12'b000000000000;
font0[1020] = 12'b000000000000;
font0[1021] = 12'b000000000000;
font0[1022] = 12'b000000000000;
font0[1023] = 12'b000000000000;
font0[1024] = 12'b000000000000;
font0[1025] = 12'b000000000000;
font0[1026] = 12'b000100001000;
font0[1027] = 12'b000100001000;
font0[1028] = 12'b000100001000;
font0[1029] = 12'b000000001000;
font0[1030] = 12'b000011111000;
font0[1031] = 12'b000000011000;
font0[1032] = 12'b000000011000;
font0[1033] = 12'b000011110000;
font0[1034] = 12'b000000000000;
font0[1035] = 12'b000000000000;
font0[1036] = 12'b000000000000;
font0[1037] = 12'b000000000000;
font0[1038] = 12'b000000000000;
font0[1039] = 12'b000000000000;
font0[1040] = 12'b000000000000;
font0[1041] = 12'b000000000000;
font0[1042] = 12'b000000000000;
font0[1043] = 12'b000000000000;
font0[1044] = 12'b001111111000;
font0[1045] = 12'b000000111000;
font0[1046] = 12'b000000110000;
font0[1047] = 12'b000001100000;
font0[1048] = 12'b000110000000;
font0[1049] = 12'b000100000000;
font0[1050] = 12'b001100000000;
font0[1051] = 12'b001111111000;
font0[1052] = 12'b000000000000;
font0[1053] = 12'b000000000000;
font0[1054] = 12'b000000000000;
font0[1055] = 12'b000000000000;
font0[1056] = 12'b000000000000;
font0[1057] = 12'b000000000000;
font0[1058] = 12'b000000000000;
font0[1059] = 12'b000000000000;
font0[1060] = 12'b000000000000;
font0[1061] = 12'b000000000000;
font0[1062] = 12'b000011110000;
font0[1063] = 12'b000010000000;
font0[1064] = 12'b000010000000;
font0[1065] = 12'b000011000000;
font0[1066] = 12'b000011000000;
font0[1067] = 12'b000011000000;
font0[1068] = 12'b000011000000;
font0[1069] = 12'b000011110000;
font0[1070] = 12'b000000000000;
font0[1071] = 12'b000000000000;
font0[1072] = 12'b000000000000;
font0[1073] = 12'b000000000000;
font0[1074] = 12'b000000000000;
font0[1075] = 12'b000000000000;
font0[1076] = 12'b000000000000;
font0[1077] = 12'b000000000000;
font0[1078] = 12'b000000000000;
font0[1079] = 12'b000000000000;
font0[1080] = 12'b000000000000;
font0[1081] = 12'b000010000000;
font0[1082] = 12'b000010000000;
font0[1083] = 12'b000001000000;
font0[1084] = 12'b000001100000;
font0[1085] = 12'b000001100000;
font0[1086] = 12'b000000110000;
font0[1087] = 12'b000000110000;
font0[1088] = 12'b000000000000;
font0[1089] = 12'b000000000000;
font0[1090] = 12'b000000000000;
font0[1091] = 12'b000000000000;
font0[1092] = 12'b000000000000;
font0[1093] = 12'b000000000000;
font0[1094] = 12'b000000000000;
font0[1095] = 12'b000000000000;
font0[1096] = 12'b000000000000;
font0[1097] = 12'b000000000000;
font0[1098] = 12'b000011110000;
font0[1099] = 12'b000000010000;
font0[1100] = 12'b000000010000;
font0[1101] = 12'b000000110000;
font0[1102] = 12'b000000110000;
font0[1103] = 12'b000000110000;
font0[1104] = 12'b000000110000;
font0[1105] = 12'b000011110000;
font0[1106] = 12'b000000000000;
font0[1107] = 12'b000000000000;
font0[1108] = 12'b000000000000;
font0[1109] = 12'b000000000000;
font0[1110] = 12'b000000000000;
font0[1111] = 12'b000000000000;
font0[1112] = 12'b000000000000;
font0[1113] = 12'b000000000000;
font0[1114] = 12'b000000000000;
font0[1115] = 12'b000000000000;
font0[1116] = 12'b000011000000;
font0[1117] = 12'b000111100000;
font0[1118] = 12'b001100110000;
font0[1119] = 12'b001000011000;
font0[1120] = 12'b000000000000;
font0[1121] = 12'b000000000000;
font0[1122] = 12'b000000000000;
font0[1123] = 12'b000000000000;
font0[1124] = 12'b000000000000;
font0[1125] = 12'b000000000000;
font0[1126] = 12'b000000000000;
font0[1127] = 12'b000000000000;
font0[1128] = 12'b000000000000;
font0[1129] = 12'b000000000000;
font0[1130] = 12'b000000000000;
font0[1131] = 12'b000000000000;
font0[1132] = 12'b000000000000;
font0[1133] = 12'b000000000000;
font0[1134] = 12'b000000000000;
font0[1135] = 12'b000000000000;
font0[1136] = 12'b000000000000;
font0[1137] = 12'b000000000000;
font0[1138] = 12'b000000000000;
font0[1139] = 12'b000000000000;
font0[1140] = 12'b000000000000;
font0[1141] = 12'b001111111000;
font0[1142] = 12'b000000000000;
font0[1143] = 12'b000000000000;
font0[1144] = 12'b000000000000;
font0[1145] = 12'b000000000000;
font0[1146] = 12'b000000000000;
font0[1147] = 12'b000000000000;
font0[1148] = 12'b000000000000;
font0[1149] = 12'b000000000000;
font0[1150] = 12'b000000000000;
font0[1151] = 12'b000000000000;
font0[1152] = 12'b000010000000;
font0[1153] = 12'b000011000000;
font0[1154] = 12'b000001100000;
font0[1155] = 12'b000000000000;
font0[1156] = 12'b000000000000;
font0[1157] = 12'b000000000000;
font0[1158] = 12'b000000000000;
font0[1159] = 12'b000000000000;
font0[1160] = 12'b000000000000;
font0[1161] = 12'b000000000000;
font0[1162] = 12'b000000000000;
font0[1163] = 12'b000000000000;
font0[1164] = 12'b000000000000;
font0[1165] = 12'b000000000000;
font0[1166] = 12'b000000000000;
font0[1167] = 12'b000000000000;
font0[1168] = 12'b000000000000;
font0[1169] = 12'b000000000000;
font0[1170] = 12'b000000000000;
font0[1171] = 12'b000000000000;
font0[1172] = 12'b000011111000;
font0[1173] = 12'b000000011000;
font0[1174] = 12'b000111111000;
font0[1175] = 12'b000100111000;
font0[1176] = 12'b000100111000;
font0[1177] = 12'b000011111000;
font0[1178] = 12'b000000000000;
font0[1179] = 12'b000000000000;
font0[1180] = 12'b000000000000;
font0[1181] = 12'b000000000000;
font0[1182] = 12'b000000000000;
font0[1183] = 12'b000000000000;
font0[1184] = 12'b000000000000;
font0[1185] = 12'b000000000000;
font0[1186] = 12'b000000000000;
font0[1187] = 12'b000000000000;
font0[1188] = 12'b000100000000;
font0[1189] = 12'b000100000000;
font0[1190] = 12'b000111110000;
font0[1191] = 12'b000110001000;
font0[1192] = 12'b000110001000;
font0[1193] = 12'b000110001000;
font0[1194] = 12'b000110001000;
font0[1195] = 12'b000111110000;
font0[1196] = 12'b000000000000;
font0[1197] = 12'b000000000000;
font0[1198] = 12'b000000000000;
font0[1199] = 12'b000000000000;
font0[1200] = 12'b000000000000;
font0[1201] = 12'b000000000000;
font0[1202] = 12'b000000000000;
font0[1203] = 12'b000000000000;
font0[1204] = 12'b000000000000;
font0[1205] = 12'b000000000000;
font0[1206] = 12'b000000000000;
font0[1207] = 12'b000000000000;
font0[1208] = 12'b000011111000;
font0[1209] = 12'b000110000000;
font0[1210] = 12'b000110000000;
font0[1211] = 12'b000110000000;
font0[1212] = 12'b000110000000;
font0[1213] = 12'b000011111000;
font0[1214] = 12'b000000000000;
font0[1215] = 12'b000000000000;
font0[1216] = 12'b000000000000;
font0[1217] = 12'b000000000000;
font0[1218] = 12'b000000000000;
font0[1219] = 12'b000000000000;
font0[1220] = 12'b000000000000;
font0[1221] = 12'b000000000000;
font0[1222] = 12'b000000000000;
font0[1223] = 12'b000000000000;
font0[1224] = 12'b000000001000;
font0[1225] = 12'b000000001000;
font0[1226] = 12'b000011111000;
font0[1227] = 12'b000100011000;
font0[1228] = 12'b000100011000;
font0[1229] = 12'b000100011000;
font0[1230] = 12'b000100011000;
font0[1231] = 12'b000011111000;
font0[1232] = 12'b000000000000;
font0[1233] = 12'b000000000000;
font0[1234] = 12'b000000000000;
font0[1235] = 12'b000000000000;
font0[1236] = 12'b000000000000;
font0[1237] = 12'b000000000000;
font0[1238] = 12'b000000000000;
font0[1239] = 12'b000000000000;
font0[1240] = 12'b000000000000;
font0[1241] = 12'b000000000000;
font0[1242] = 12'b000000000000;
font0[1243] = 12'b000000000000;
font0[1244] = 12'b000011110000;
font0[1245] = 12'b000111001000;
font0[1246] = 12'b000111001000;
font0[1247] = 12'b000111111000;
font0[1248] = 12'b000111000000;
font0[1249] = 12'b000011110000;
font0[1250] = 12'b000000000000;
font0[1251] = 12'b000000000000;
font0[1252] = 12'b000000000000;
font0[1253] = 12'b000000000000;
font0[1254] = 12'b000000000000;
font0[1255] = 12'b000000000000;
font0[1256] = 12'b000000000000;
font0[1257] = 12'b000000000000;
font0[1258] = 12'b000000000000;
font0[1259] = 12'b000000000000;
font0[1260] = 12'b000001110000;
font0[1261] = 12'b000010011000;
font0[1262] = 12'b000010000000;
font0[1263] = 12'b000010000000;
font0[1264] = 12'b000111110000;
font0[1265] = 12'b000011000000;
font0[1266] = 12'b000011000000;
font0[1267] = 12'b000011000000;
font0[1268] = 12'b000000000000;
font0[1269] = 12'b000000000000;
font0[1270] = 12'b000000000000;
font0[1271] = 12'b000000000000;
font0[1272] = 12'b000000000000;
font0[1273] = 12'b000000000000;
font0[1274] = 12'b000000000000;
font0[1275] = 12'b000000000000;
font0[1276] = 12'b000000000000;
font0[1277] = 12'b000000000000;
font0[1278] = 12'b000000000000;
font0[1279] = 12'b000000000000;
font0[1280] = 12'b000011110000;
font0[1281] = 12'b000100111000;
font0[1282] = 12'b000100111000;
font0[1283] = 12'b000100111000;
font0[1284] = 12'b000100111000;
font0[1285] = 12'b000011111000;
font0[1286] = 12'b000000111000;
font0[1287] = 12'b000011110000;
font0[1288] = 12'b000000000000;
font0[1289] = 12'b000000000000;
font0[1290] = 12'b000000000000;
font0[1291] = 12'b000000000000;
font0[1292] = 12'b000000000000;
font0[1293] = 12'b000000000000;
font0[1294] = 12'b000000000000;
font0[1295] = 12'b000000000000;
font0[1296] = 12'b000100000000;
font0[1297] = 12'b000100000000;
font0[1298] = 12'b000111110000;
font0[1299] = 12'b000100001000;
font0[1300] = 12'b000110001000;
font0[1301] = 12'b000110001000;
font0[1302] = 12'b000110001000;
font0[1303] = 12'b000110001000;
font0[1304] = 12'b000000000000;
font0[1305] = 12'b000000000000;
font0[1306] = 12'b000000000000;
font0[1307] = 12'b000000000000;
font0[1308] = 12'b000000000000;
font0[1309] = 12'b000000000000;
font0[1310] = 12'b000000000000;
font0[1311] = 12'b000000000000;
font0[1312] = 12'b000000000000;
font0[1313] = 12'b000000000000;
font0[1314] = 12'b000001100000;
font0[1315] = 12'b000000000000;
font0[1316] = 12'b000011110000;
font0[1317] = 12'b000001100000;
font0[1318] = 12'b000001100000;
font0[1319] = 12'b000001100000;
font0[1320] = 12'b000001100000;
font0[1321] = 12'b000011110000;
font0[1322] = 12'b000000000000;
font0[1323] = 12'b000000000000;
font0[1324] = 12'b000000000000;
font0[1325] = 12'b000000000000;
font0[1326] = 12'b000000000000;
font0[1327] = 12'b000000000000;
font0[1328] = 12'b000000000000;
font0[1329] = 12'b000000000000;
font0[1330] = 12'b000000000000;
font0[1331] = 12'b000000000000;
font0[1332] = 12'b000001100000;
font0[1333] = 12'b000000000000;
font0[1334] = 12'b000011110000;
font0[1335] = 12'b000000110000;
font0[1336] = 12'b000000110000;
font0[1337] = 12'b000000110000;
font0[1338] = 12'b000000110000;
font0[1339] = 12'b000000110000;
font0[1340] = 12'b000110110000;
font0[1341] = 12'b000011100000;
font0[1342] = 12'b000000000000;
font0[1343] = 12'b000000000000;
font0[1344] = 12'b000000000000;
font0[1345] = 12'b000000000000;
font0[1346] = 12'b000000000000;
font0[1347] = 12'b000000000000;
font0[1348] = 12'b000000000000;
font0[1349] = 12'b000000000000;
font0[1350] = 12'b000100000000;
font0[1351] = 12'b000100000000;
font0[1352] = 12'b000100001000;
font0[1353] = 12'b000100001000;
font0[1354] = 12'b000111100000;
font0[1355] = 12'b000110010000;
font0[1356] = 12'b000110001000;
font0[1357] = 12'b000110001000;
font0[1358] = 12'b000000000000;
font0[1359] = 12'b000000000000;
font0[1360] = 12'b000000000000;
font0[1361] = 12'b000000000000;
font0[1362] = 12'b000000000000;
font0[1363] = 12'b000000000000;
font0[1364] = 12'b000000000000;
font0[1365] = 12'b000000000000;
font0[1366] = 12'b000000000000;
font0[1367] = 12'b000000000000;
font0[1368] = 12'b000011000000;
font0[1369] = 12'b000001000000;
font0[1370] = 12'b000001000000;
font0[1371] = 12'b000001100000;
font0[1372] = 12'b000001100000;
font0[1373] = 12'b000001100000;
font0[1374] = 12'b000001100000;
font0[1375] = 12'b000011110000;
font0[1376] = 12'b000000000000;
font0[1377] = 12'b000000000000;
font0[1378] = 12'b000000000000;
font0[1379] = 12'b000000000000;
font0[1380] = 12'b000000000000;
font0[1381] = 12'b000000000000;
font0[1382] = 12'b000000000000;
font0[1383] = 12'b000000000000;
font0[1384] = 12'b000000000000;
font0[1385] = 12'b000000000000;
font0[1386] = 12'b000000000000;
font0[1387] = 12'b000000000000;
font0[1388] = 12'b001111111000;
font0[1389] = 12'b001100100100;
font0[1390] = 12'b001110100100;
font0[1391] = 12'b001110100100;
font0[1392] = 12'b001110100100;
font0[1393] = 12'b001110100100;
font0[1394] = 12'b000000000000;
font0[1395] = 12'b000000000000;
font0[1396] = 12'b000000000000;
font0[1397] = 12'b000000000000;
font0[1398] = 12'b000000000000;
font0[1399] = 12'b000000000000;
font0[1400] = 12'b000000000000;
font0[1401] = 12'b000000000000;
font0[1402] = 12'b000000000000;
font0[1403] = 12'b000000000000;
font0[1404] = 12'b000000000000;
font0[1405] = 12'b000000000000;
font0[1406] = 12'b000111110000;
font0[1407] = 12'b000110001000;
font0[1408] = 12'b000111001000;
font0[1409] = 12'b000111001000;
font0[1410] = 12'b000111001000;
font0[1411] = 12'b000111001000;
font0[1412] = 12'b000000000000;
font0[1413] = 12'b000000000000;
font0[1414] = 12'b000000000000;
font0[1415] = 12'b000000000000;
font0[1416] = 12'b000000000000;
font0[1417] = 12'b000000000000;
font0[1418] = 12'b000000000000;
font0[1419] = 12'b000000000000;
font0[1420] = 12'b000000000000;
font0[1421] = 12'b000000000000;
font0[1422] = 12'b000000000000;
font0[1423] = 12'b000000000000;
font0[1424] = 12'b000011110000;
font0[1425] = 12'b000111001000;
font0[1426] = 12'b000111001000;
font0[1427] = 12'b000111001000;
font0[1428] = 12'b000111001000;
font0[1429] = 12'b000011110000;
font0[1430] = 12'b000000000000;
font0[1431] = 12'b000000000000;
font0[1432] = 12'b000000000000;
font0[1433] = 12'b000000000000;
font0[1434] = 12'b000000000000;
font0[1435] = 12'b000000000000;
font0[1436] = 12'b000000000000;
font0[1437] = 12'b000000000000;
font0[1438] = 12'b000000000000;
font0[1439] = 12'b000000000000;
font0[1440] = 12'b000000000000;
font0[1441] = 12'b000000000000;
font0[1442] = 12'b000111110000;
font0[1443] = 12'b000110001000;
font0[1444] = 12'b000111001000;
font0[1445] = 12'b000111001000;
font0[1446] = 12'b000111001000;
font0[1447] = 12'b000111110000;
font0[1448] = 12'b000111000000;
font0[1449] = 12'b000111000000;
font0[1450] = 12'b000000000000;
font0[1451] = 12'b000000000000;
font0[1452] = 12'b000000000000;
font0[1453] = 12'b000000000000;
font0[1454] = 12'b000000000000;
font0[1455] = 12'b000000000000;
font0[1456] = 12'b000000000000;
font0[1457] = 12'b000000000000;
font0[1458] = 12'b000000000000;
font0[1459] = 12'b000000000000;
font0[1460] = 12'b000011111000;
font0[1461] = 12'b000100011000;
font0[1462] = 12'b000100111000;
font0[1463] = 12'b000100111000;
font0[1464] = 12'b000100111000;
font0[1465] = 12'b000011111000;
font0[1466] = 12'b000000111000;
font0[1467] = 12'b000000111000;
font0[1468] = 12'b000000000000;
font0[1469] = 12'b000000000000;
font0[1470] = 12'b000000000000;
font0[1471] = 12'b000000000000;
font0[1472] = 12'b000000000000;
font0[1473] = 12'b000000000000;
font0[1474] = 12'b000000000000;
font0[1475] = 12'b000000000000;
font0[1476] = 12'b000000000000;
font0[1477] = 12'b000000000000;
font0[1478] = 12'b000111110000;
font0[1479] = 12'b000100011000;
font0[1480] = 12'b000110000000;
font0[1481] = 12'b000110000000;
font0[1482] = 12'b000110000000;
font0[1483] = 12'b000110000000;
font0[1484] = 12'b000000000000;
font0[1485] = 12'b000000000000;
font0[1486] = 12'b000000000000;
font0[1487] = 12'b000000000000;
font0[1488] = 12'b000000000000;
font0[1489] = 12'b000000000000;
font0[1490] = 12'b000000000000;
font0[1491] = 12'b000000000000;
font0[1492] = 12'b000000000000;
font0[1493] = 12'b000000000000;
font0[1494] = 12'b000000000000;
font0[1495] = 12'b000000000000;
font0[1496] = 12'b000011111000;
font0[1497] = 12'b000100000000;
font0[1498] = 12'b000111110000;
font0[1499] = 12'b000000011000;
font0[1500] = 12'b000000011000;
font0[1501] = 12'b000111110000;
font0[1502] = 12'b000000000000;
font0[1503] = 12'b000000000000;
font0[1504] = 12'b000000000000;
font0[1505] = 12'b000000000000;
font0[1506] = 12'b000000000000;
font0[1507] = 12'b000000000000;
font0[1508] = 12'b000000000000;
font0[1509] = 12'b000000000000;
font0[1510] = 12'b000000000000;
font0[1511] = 12'b000000000000;
font0[1512] = 12'b000010000000;
font0[1513] = 12'b000010000000;
font0[1514] = 12'b000010000000;
font0[1515] = 12'b000111110000;
font0[1516] = 12'b000011000000;
font0[1517] = 12'b000011000000;
font0[1518] = 12'b000011011000;
font0[1519] = 12'b000001110000;
font0[1520] = 12'b000000000000;
font0[1521] = 12'b000000000000;
font0[1522] = 12'b000000000000;
font0[1523] = 12'b000000000000;
font0[1524] = 12'b000000000000;
font0[1525] = 12'b000000000000;
font0[1526] = 12'b000000000000;
font0[1527] = 12'b000000000000;
font0[1528] = 12'b000000000000;
font0[1529] = 12'b000000000000;
font0[1530] = 12'b000000000000;
font0[1531] = 12'b000000000000;
font0[1532] = 12'b000110001000;
font0[1533] = 12'b000111001000;
font0[1534] = 12'b000111001000;
font0[1535] = 12'b000111001000;
font0[1536] = 12'b000111001000;
font0[1537] = 12'b000011110000;
font0[1538] = 12'b000000000000;
font0[1539] = 12'b000000000000;
font0[1540] = 12'b000000000000;
font0[1541] = 12'b000000000000;
font0[1542] = 12'b000000000000;
font0[1543] = 12'b000000000000;
font0[1544] = 12'b000000000000;
font0[1545] = 12'b000000000000;
font0[1546] = 12'b000000000000;
font0[1547] = 12'b000000000000;
font0[1548] = 12'b000000000000;
font0[1549] = 12'b000000000000;
font0[1550] = 12'b000110001000;
font0[1551] = 12'b000111001000;
font0[1552] = 12'b000111001000;
font0[1553] = 12'b000111001000;
font0[1554] = 12'b000011010000;
font0[1555] = 12'b000001110000;
font0[1556] = 12'b000000000000;
font0[1557] = 12'b000000000000;
font0[1558] = 12'b000000000000;
font0[1559] = 12'b000000000000;
font0[1560] = 12'b000000000000;
font0[1561] = 12'b000000000000;
font0[1562] = 12'b000000000000;
font0[1563] = 12'b000000000000;
font0[1564] = 12'b000000000000;
font0[1565] = 12'b000000000000;
font0[1566] = 12'b000000000000;
font0[1567] = 12'b000000000000;
font0[1568] = 12'b001100000100;
font0[1569] = 12'b001110100100;
font0[1570] = 12'b001110100100;
font0[1571] = 12'b001110100100;
font0[1572] = 12'b001110100100;
font0[1573] = 12'b000111111000;
font0[1574] = 12'b000000000000;
font0[1575] = 12'b000000000000;
font0[1576] = 12'b000000000000;
font0[1577] = 12'b000000000000;
font0[1578] = 12'b000000000000;
font0[1579] = 12'b000000000000;
font0[1580] = 12'b000000000000;
font0[1581] = 12'b000000000000;
font0[1582] = 12'b000000000000;
font0[1583] = 12'b000000000000;
font0[1584] = 12'b000000000000;
font0[1585] = 12'b000000000000;
font0[1586] = 12'b000110111000;
font0[1587] = 12'b000110111000;
font0[1588] = 12'b000011100000;
font0[1589] = 12'b000010110000;
font0[1590] = 12'b000110111000;
font0[1591] = 12'b000110111000;
font0[1592] = 12'b000000000000;
font0[1593] = 12'b000000000000;
font0[1594] = 12'b000000000000;
font0[1595] = 12'b000000000000;
font0[1596] = 12'b000000000000;
font0[1597] = 12'b000000000000;
font0[1598] = 12'b000000000000;
font0[1599] = 12'b000000000000;
font0[1600] = 12'b000000000000;
font0[1601] = 12'b000000000000;
font0[1602] = 12'b000000000000;
font0[1603] = 12'b000000000000;
font0[1604] = 12'b000100111000;
font0[1605] = 12'b000100111000;
font0[1606] = 12'b000100111000;
font0[1607] = 12'b000100111000;
font0[1608] = 12'b000100111000;
font0[1609] = 12'b000011111000;
font0[1610] = 12'b000000111000;
font0[1611] = 12'b000011110000;
font0[1612] = 12'b000000000000;
font0[1613] = 12'b000000000000;
font0[1614] = 12'b000000000000;
font0[1615] = 12'b000000000000;
font0[1616] = 12'b000000000000;
font0[1617] = 12'b000000000000;
font0[1618] = 12'b000000000000;
font0[1619] = 12'b000000000000;
font0[1620] = 12'b000000000000;
font0[1621] = 12'b000000000000;
font0[1622] = 12'b000111111000;
font0[1623] = 12'b000000111000;
font0[1624] = 12'b000011100000;
font0[1625] = 12'b000010000000;
font0[1626] = 12'b000110000000;
font0[1627] = 12'b000111111000;
font0[1628] = 12'b000000000000;
font0[1629] = 12'b000000000000;
font0[1630] = 12'b000000000000;
font0[1631] = 12'b000000000000;
font0[1632] = 12'b000000000000;
font0[1633] = 12'b000000000000;
font0[1634] = 12'b000000000000;
font0[1635] = 12'b000000000000;
font0[1636] = 12'b000000000000;
font0[1637] = 12'b000000000000;
font0[1638] = 12'b000011110000;
font0[1639] = 12'b000010000000;
font0[1640] = 12'b000010000000;
font0[1641] = 12'b000010000000;
font0[1642] = 12'b000111000000;
font0[1643] = 12'b000011000000;
font0[1644] = 12'b000011000000;
font0[1645] = 12'b000011110000;
font0[1646] = 12'b000000000000;
font0[1647] = 12'b000000000000;
font0[1648] = 12'b000000000000;
font0[1649] = 12'b000000000000;
font0[1650] = 12'b000000000000;
font0[1651] = 12'b000000000000;
font0[1652] = 12'b000000000000;
font0[1653] = 12'b000000000000;
font0[1654] = 12'b000000000000;
font0[1655] = 12'b000000000000;
font0[1656] = 12'b000001000000;
font0[1657] = 12'b000001000000;
font0[1658] = 12'b000001000000;
font0[1659] = 12'b000001000000;
font0[1660] = 12'b000001100000;
font0[1661] = 12'b000001100000;
font0[1662] = 12'b000001100000;
font0[1663] = 12'b000001100000;
font0[1664] = 12'b000000000000;
font0[1665] = 12'b000000000000;
font0[1666] = 12'b000000000000;
font0[1667] = 12'b000000000000;
font0[1668] = 12'b000000000000;
font0[1669] = 12'b000000000000;
font0[1670] = 12'b000000000000;
font0[1671] = 12'b000000000000;
font0[1672] = 12'b000000000000;
font0[1673] = 12'b000000000000;
font0[1674] = 12'b000111100000;
font0[1675] = 12'b000000100000;
font0[1676] = 12'b000000100000;
font0[1677] = 12'b000000100000;
font0[1678] = 12'b000001110000;
font0[1679] = 12'b000001100000;
font0[1680] = 12'b000001100000;
font0[1681] = 12'b000111100000;
font0[1682] = 12'b000000000000;
font0[1683] = 12'b000000000000;
font0[1684] = 12'b000000000000;
font0[1685] = 12'b000000000000;
font0[1686] = 12'b000000000000;
font0[1687] = 12'b000000000000;
font0[1688] = 12'b000000000000;
font0[1689] = 12'b000000000000;
font0[1690] = 12'b000000000000;
font0[1691] = 12'b000000000000;
font0[1692] = 12'b000000000000;
font0[1693] = 12'b000000000000;
font0[1694] = 12'b000110000000;
font0[1695] = 12'b001001001000;
font0[1696] = 12'b001001111000;
font0[1697] = 12'b000000000000;
font0[1698] = 12'b000000000000;
font0[1699] = 12'b000000000000;
font0[1700] = 12'b000000000000;
font0[1701] = 12'b000000000000;
font0[1702] = 12'b000000000000;
font0[1703] = 12'b000000000000;
font0[1704] = 12'b000000000000;
font0[1705] = 12'b000000000000;
font0[1706] = 12'b000000000000;
font0[1707] = 12'b000000000000;
font0[1708] = 12'b000000000000;
font0[1709] = 12'b000000000000;
end
/* #### END FONT0 #### */
