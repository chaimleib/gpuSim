`define GPU_Swap            (1)
`define GPU_ChangeColorMap  (0)
`define GPU_Pixel           (2)
`define GPU_Rect            (3)

