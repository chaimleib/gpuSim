`define TestVectorCount (580)

